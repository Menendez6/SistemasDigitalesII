



suma1 = signed(ent_a(7 downto 0)) + signed (ent_b(7 downto 0));

suma <= "01111111" when suma1(7) = '1'